package constants is

	-- delay for logic gates
	constant IVDELAY : time := 0.1 ns;
	constant NDDELAY : time := 0.2 ns;
	
	-- default number of bits
	constant Nbit : integer := 4;
	
end constants;