package constants is

	-- delay for logic gates
	constant IVDELAY : time := 0.1 ns;
	constant NDDELAY : time := 0.2 ns;
	
	-- default number of bits
	constant numBit : integer := 4;

	-- delay mux
	constant tp_mux : time := 0.5 ns;
	
end constants;
